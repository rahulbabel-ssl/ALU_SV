package alu_package;
        `include "alu_transaction.sv"
        `include "alu_generator.sv"
        `include "alu_monitor.sv"
        `include "alu_driver.sv"
        `include "alu_scoreboard.sv"
        `include "alu_reference.sv"
        `include "alu_environment.sv"
        `include "alu_test.sv"
        endpackage
